LIBRARY IEEE;
LIBRARY work;
USE IEEE.fixed_float_types.ALL;
USE IEEE.fixed_pkg.ALL;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE IEEE.std_logic_unsigned.ALL;
USE work.c_pkg.ALL;

ENTITY pool_window IS
	GENERIC (FILTER_SIZE : INTEGER := 2;IMG_SIZE : INTEGER := 4);
	PORT(
		IMG :  IN STD_LOGIC_VECTOR((IMG_SIZE*IMG_SIZE*16)-1 DOWNTO 0);
		clk , START , rst :IN STD_LOGIC;
		Done : OUT STD_LOGIC;
		pool_img : OUT STD_LOGIC_VECTOR((IMG_SIZE/2)*(IMG_SIZE/2)*16-1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE pool_image_arch OF pool_window IS

	COMPONENT extract_window IS
		GENERIC (FILTER_SIZE : INTEGER ;IMG_SIZE : INTEGER);
		PORT(
			IMG : IN STD_LOGIC_VECTOR(IMG_SIZE*IMG_SIZE*16-1 DOWNTO 0);
			IMG_SIZE_in:IN INTEGER;
			FILTER_SIZE_in:IN INTEGER;
			rst:IN STD_LOGIC;
			OFFSET:IN INTEGER;
			LAYER : OUT STD_LOGIC_VECTOR(FILTER_SIZE*FILTER_SIZE*16-1 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT Pool IS
		GENERIC (WINDOW_SIZE : INTEGER := 2);
		PORT(
			WINDOW : IN STD_LOGIC_VECTOR((WINDOW_SIZE*WINDOW_SIZE*16)-1 DOWNTO 0);
			START,rst,clk : IN STD_LOGIC;
			AVR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			Done : OUT STD_LOGIC
		);
	END COMPONENT;

	TYPE conv_type IS ARRAY(0 TO ((IMG_SIZE/2)*(IMG_SIZE/2) -1))OF STD_LOGIC_VECTOR(FILTER_SIZE*FILTER_SIZE*16-1 DOWNTO 0);
	TYPE OFFSSET_type IS ARRAY(0 TO ((IMG_SIZE/2)*(IMG_SIZE/2) -1)) OF unsigned(9 DOWNTO 0);

	SIGNAL WINDOW : conv_type;
	SIGNAL OFFSSET : OFFSSET_type ;
	SIGNAL MiniPoolDone,temp1 : STD_LOGIC_VECTOR(0 TO (IMG_SIZE/2)*(IMG_SIZE/2)-1);
		
	BEGIN
		OFFSSET(0)<=(OTHERS =>'0');	
		loop0: FOR i IN 1 TO (IMG_SIZE/2)*(IMG_SIZE/2)-1 GENERATE 
			OFFSSET(i) <= OFFSSET(i-1)+"0000000010"+IMG_SIZE when( (to_integer(OFFSSET(i-1))+FILTER_SIZE )mod  IMG_SIZE)=0 ELSE
			OFFSSET(i-1)+"0000000010" ;
		END GENERATE;

		loop1: FOR i IN 0 TO (IMG_SIZE/2)*(IMG_SIZE/2)-1  GENERATE 
			fx0:extract_window GENERIC MAP (FILTER_SIZE,IMG_SIZE)PORT MAP(IMG,IMG_SIZE,FILTER_SIZE,rst,to_integer(OFFSSET(i)),WINDOW(i));

			fx1:Pool GENERIC MAP (FILTER_SIZE) PORT MAP(WINDOW(i),START,rst,clk,pool_img(i*16+15 DOWNTO i*16),MiniPoolDone(i));

		END GENERATE;

		temp1 <= (OTHERS => '1');
		Done <= '1' WHEN MiniPoolDone = temp1
				  ELSE '0';

	END pool_image_arch;