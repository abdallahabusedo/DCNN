LIBRARY IEEE;
LIBRARY work;
USE IEEE.fixed_float_types.ALL;
USE IEEE.fixed_pkg.ALL;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE IEEE.std_logic_unsigned.ALL;

ENTITY convolut_image IS
GENERIC (FILTER_SIZE : INTEGER := 3;IMG_SIZE : INTEGER := 5);
	PORT(
		IMG : IN  STD_LOGIC_VECTOR(IMG_SIZE*IMG_SIZE*16-1 DOWNTO 0);
		FILTER1 : IN STD_LOGIC_VECTOR(FILTER_SIZE*FILTER_SIZE*16-1 DOWNTO 0);
		convoluted_img : OUT STD_LOGIC_VECTOR((IMG_SIZE-FILTER_SIZE+1)*(IMG_SIZE-FILTER_SIZE+1)*16-1 DOWNTO 0);
		end_conv :OUT STD_LOGIC;
		clk,strat_signal,REST:IN STD_LOGIC
	);
END ENTITY;
ARCHITECTURE conv_image_arch OF convolut_image IS
COMPONENT conv_wimdow_1 IS 
	GENERIC (FILTER_SIZE : INTEGER);
	PORT(
		WINDOW : IN STD_LOGIC_VECTOR(FILTER_SIZE*FILTER_SIZE*16-1 DOWNTO 0);
		FILTER : IN STD_LOGIC_VECTOR(FILTER_SIZE*FILTER_SIZE*16-1 DOWNTO 0);
		PIXEL_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		end_conv :OUT STD_LOGIC;
		clk,strat_signal,REST:IN STD_LOGIC
	);
END COMPONENT;
----------------------------------------------------
COMPONENT extract_window IS
	PORT(
		IMG : IN STD_LOGIC_VECTOR(IMG_SIZE*IMG_SIZE*16-1 DOWNTO 0);
		IMG_SIZE_in:IN INTEGER;
		FILTER_SIZE_in:IN INTEGER;
		REST:IN STD_LOGIC;
		OFFSET:IN INTEGER;
		LAYER : OUT STD_LOGIC_VECTOR(FILTER_SIZE*FILTER_SIZE*16-1 DOWNTO 0)
	);
END COMPONENT;

TYPE conv_type IS ARRAY(0 TO (IMG_SIZE-FILTER_SIZE+1)*(IMG_SIZE-FILTER_SIZE+1)-1)OF STD_LOGIC_VECTOR(FILTER_SIZE*FILTER_SIZE*16-1 DOWNTO 0);
SIGNAL WINDOW : conv_type;
SIGNAL y: STD_LOGIC_VECTOR((IMG_SIZE-FILTER_SIZE+1)*(IMG_SIZE-FILTER_SIZE+1)*16-1 DOWNTO 0);

TYPE OFFSSET_type IS ARRAY(0 TO (IMG_SIZE-FILTER_SIZE+1)*(IMG_SIZE-FILTER_SIZE+1)-1) OF unsigned(9 DOWNTO 0);
	SIGNAL OFFSSET : OFFSSET_type ;
	BEGIN
		OFFSSET(0)<=(OTHERS =>'0');	
		loop0: FOR i IN 1 TO (IMG_SIZE-FILTER_SIZE+1)*(IMG_SIZE-FILTER_SIZE+1)-1 GENERATE 		
				OFFSSET(i) <= OFFSSET(i-1)+to_unsigned(FILTER_SIZE,10) WHEN ( (to_integer(OFFSSET(i-1))+FILTER_SIZE )mod  IMG_SIZE)=0 else
       				OFFSSET(i-1)+"0000000001" ;
		END GENERATE;
		loop1: FOR i IN 0 TO (IMG_SIZE-FILTER_SIZE+1)*(IMG_SIZE-FILTER_SIZE+1)-1   GENERATE 		
				fx0:extract_window GENERIC MAP (FILTER_SIZE,IMG_SIZE)PORT MAP(IMG,IMG_SIZE,FILTER_SIZE,REST,to_integer(OFFSSET(i)),WINDOW(i));
				fx1:conv_wimdow_1 GENERIC MAP (FILTER_SIZE)  PORT MAP(WINDOW(i),
					FILTER1,convoluted_img(i*16+15 DOWNTO i*16),end_conv,clk,strat_signal,REST);
   	
		END GENERATE;
END conv_image_arch;

